`define Enable        1'b1
`define Disable       1'b0
`define ZeroWord      32'b0   // 默认的零信息
`define ZeroByte      8'b0 